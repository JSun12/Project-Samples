module flash_fsm (clk, pause, play_forward, restart, sync_clk_edge, waitrequest, data_valid, flash_data, read, read_address, audio_data, kbd_rst, interrupt_event);
input clk;   //clock the fsm will run at
input pause;    //whether or not to pause music play back
input play_forward;   //whether or not to play in reverse
input restart;    //whether or not to restart song
input sync_clk_edge;    //rising edge of the clock the music will play at
input waitrequest;    //wait request generated by flash memory module
input data_valid;   //data validity flag generated by flash memory module
input [31:0] flash_data;    //data read from flash memory
output reg read;    //read flag for the flash memory to use
output reg [22:0] read_address;   //address in the flash memory to read from
output reg [7:0] audio_data;    //digital data to be generated to sound
output reg kbd_rst;   //flag to reset keyboard ascii data
output reg interrupt_event;
reg [6:0] state;
initial interrupt_event = 0;

//define all possible fsm states in one-hot
parameter [6:0] ASSERT      = 7'b0000001;
parameter [6:0] READ        = 7'b0000010;
parameter [6:0] PLAY_LOWER  = 7'b0000100;
parameter [6:0] DIS_ISR_1   = 7'b0001000;
parameter [6:0] PLAY_UPPER  = 7'b0010000;
parameter [6:0] DIS_ISR_2   = 7'b0100000;
parameter [6:0] UPDATE_ADDR = 7'b1000000;

//define the start and end address of the song
parameter [22:0] max_address = 23'b00001111111111111111111;
parameter [22:0] min_address = 23'b0;

//reg [4:0] state;
reg [22:0] address_counter;   //address to be incremented
initial address_counter = 23'b0;    //initialize address_counter to starting address
reg [31:0] song_data;   //data read from fsm

// assert address and read signal at clock cycle
// waitrequest -> wait for readdatavalid
// While waiting, address, read, write, and byteenable can't change
// look at readdata
always_ff @(posedge clk or posedge pause) begin
  //loop assert state if pause is high (asynchronous)
  if (pause)
    state <= ASSERT;
  else begin
  case(state)
    ASSERT:      begin
                  //set read to 1 and set read_address to incremented address
                 read <= 1'b1;
                 read_address <= address_counter;
                  //loop assert state if waitrequest is generated
                 if (waitrequest) 
                  state <= ASSERT;
                 else
                  state <= READ;
                 end
    READ:        //read data from flash memory and set read to 0 if data is valid
                 if (data_valid) begin
                   song_data <= flash_data;
                   read <= 1'b0;
                   state <= PLAY_LOWER;
                 end
                 else
                   state <= READ;
    PLAY_LOWER:  //play most significant 8 bits of the lower 16 bit flash data on posedge song clock
                 if (sync_clk_edge) begin
                   audio_data <= song_data[15:8];
                   interrupt_event <= 1'b1;       //generate interrupt event flag
                   state <= DIS_ISR_1;
                 end
                 else
                   state <= PLAY_LOWER;
    DIS_ISR_1:   begin
                   interrupt_event <= 1'b0;       //disable interrupt event flag
                   state <= PLAY_UPPER;
                 end
    PLAY_UPPER:  //play least significant 8 bits of the lower 16 bit flash data on posedge song clock
                 if (sync_clk_edge) begin
                   audio_data <= song_data[31:24];
                   interrupt_event <= 1'b1;       //generate interrupt event flag
                   state <= DIS_ISR_2;
                 end
                 else
                   state <= PLAY_UPPER;
    DIS_ISR_2:   begin
                   interrupt_event <= 1'b0;       //disable interrupt event flag
                   state <= UPDATE_ADDR;
                 end
    UPDATE_ADDR: begin
                 state <= ASSERT;
                                  //set address_counter to the starting address if restart flag is high and set kbd_rst flag to high
                 if (restart) begin
                   address_counter <= min_address;
                   kbd_rst <= 1'b1;
                 end
                 //keep going through song otherwise
                 else begin
                   kbd_rst <= 1'b0;
                 //play music forwards if play_forward flag is high
                 if (play_forward) begin
                   if (address_counter < max_address)
                     address_counter <= address_counter + 1;
                   //reset address to start at the end of the song
                   else if (address_counter >= max_address)
                     address_counter <= min_address;
                 end
                 //play music backwards if play_forward flag is low
                 else if (!play_forward) begin
                   if (address_counter > min_address)
                     address_counter <= address_counter - 1;
                   //reset address to end of the song when reversed to start
                   else if (address_counter == min_address)
                     address_counter <= max_address;
                 end
                 //this state shouldn't happen
                 else
                   address_counter <= min_address;
                 end
                 end
    default:  state <= ASSERT;
  endcase
  end
end
endmodule